//-------------------------------------------------------------------------------
//  FEUP / M.EEC - Digital Systems Design 2022/2023
//
// ADD YOUR NAMES HERE
//-------------------------------------------------------------------------------

module psddivide(
					input         clock,		//master clock
					input         reset,		//synch reset, active high
					input         start,		//start a new division
					input         stop,			//load output registers
					input  [31:0] dividend,		// dividend
					input  [31:0] divisor,		// divisor
					output [31:0] quotient,		// quotient
					output [31:0] rest			//rest
				);


// ADD YOUR CODE HERE

endmodule
